

module avalon_saber_interface (
	// Avalon Clock Input
	input logic CLK,
	// Avalon Reset Input
	input logic RESET,
	// Avalon-MM Slave Signals
	input  logic AVL_READ,					// Avalon-MM Read
	input  logic AVL_WRITE,					// Avalon-MM Write
	input  logic AVL_CS,						// Avalon-MM Chip Select
	input  logic [3:0] AVL_BYTE_EN,		// Avalon-MM Byte Enable
	input  logic [5:0] AVL_ADDR,			// Avalon-MM Address
	input  logic [31:0] AVL_WRITEDATA,	// Avalon-MM Write Data
	output logic [31:0] AVL_READDATA,	// Avalon-MM Read Data
	// Exported Conduit
	output logic [319:0] EXPORT_DATA		// Exported Conduit Signal to LEDs
);



	// create 64 32bit registers
	logic [10:0][31:0] Reg_unit;
	assign EXPORT_DATA = Reg_unit;
	always_ff @ (posedge CLK)
	begin
		if (RESET)				// if reset is active, clear all registers
			begin
				Reg_unit[0]  <= 32'h0;	// saber_exist 			  0
				Reg_unit[1]  <= 32'h0;  // saber_position x	  32
				Reg_unit[2]  <= 32'h0;  // saber_position y 	  64
				Reg_unit[3]  <= 32'h0;  // saber state			  96
				Reg_unit[4]  <= 32'h0;	// saber_figure		  128
				Reg_unit[5]  <= 32'h0;	// saber_hidden		  160
				Reg_unit[6]  <= 32'h0;	
				Reg_unit[7]  <= 32'h0;  // monster1_exist		  224
				Reg_unit[8]  <= 32'h0;  // monster1_position x 256
				Reg_unit[9]  <= 32'h0;  // monster1_position y 288
				Reg_unit[10] <= 32'h0;  // monster1_state	
			
			end

		else if (AVL_WRITE && AVL_CS)

			// Write

			begin

				case (AVL_BYTE_EN)

					4'b1111: Reg_unit[AVL_ADDR]		  <= AVL_WRITEDATA;

					4'b1100:	Reg_unit[AVL_ADDR][31:16] <= AVL_WRITEDATA[31:16];

					4'b0011: Reg_unit[AVL_ADDR][15:0]  <= AVL_WRITEDATA[15:0];

					4'b1000: Reg_unit[AVL_ADDR][31:24] <= AVL_WRITEDATA[31:24];

					4'b0100: Reg_unit[AVL_ADDR][23:16] <= AVL_WRITEDATA[23:16];

					4'b0010: Reg_unit[AVL_ADDR][15:8]  <= AVL_WRITEDATA[15:8];

					4'b0001: Reg_unit[AVL_ADDR][7:0]   <= AVL_WRITEDATA[7:0];

					default: Reg_unit[AVL_ADDR] 		  <= 32'b0;

				endcase

			end

	end

	

	

	always_comb

	begin

		AVL_READDATA = 32'b0;

		// Read

		if (AVL_READ)

			AVL_READDATA = Reg_unit[AVL_ADDR];

	end

endmodule